module encoder_1x2(
    input d0,
    input d1,
    output b
);

assign b = d1 ;

endmodule
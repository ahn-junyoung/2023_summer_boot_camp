module and (
    ports
);
    
endmodule